module D_ff_cnt( input d,output reg q);
	always@(d)
		q=d;
endmodule
